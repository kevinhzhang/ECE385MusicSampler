module ledger_line_rom (
	input [4:0] addr,
	output [7:0] data
);

	parameter ADDR_WIDTH = 5;
	parameter DATA_WIDTH = 8;
	
	parameter[0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
		  // CODE 0x00 - BLANK
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00000000, // 5
        8'b00000000, // 6
        8'b00000000, // 7
		  // CODE 0x01 - MIDDLE
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b11111111, // 4  ********
        8'b00000000, // 5
        8'b00000000, // 6
        8'b00000000, // 7 
		  // CODE 0x02 - ABOVE
        8'b11111111, // 0  ********
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00000000, // 5
        8'b00000000, // 6
        8'b00000000, // 7
		  // CODE 0x03 - BELOW
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00000000, // 5
        8'b00000000, // 6
        8'b11111111, // 7  ********
	};
	
	assign data = ROM[addr];

endmodule
