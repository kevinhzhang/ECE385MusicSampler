module note_rom (
	input [7:0] addr,
	output [7:0] data
);

	parameter ADDR_WIDTH = 5;
	parameter DATA_WIDTH = 8;
	
	// ROM definition
	parameter[0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
		  // CODE 0x00 - BLANK
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00000000, // 5
        8'b00000000, // 6
        8'b00000000, // 7
		  // CODE 0x01 - BLACK BODY ("QUARTER")
        8'b00000000, // 0
        8'b00011000, // 1     **  
        8'b01111110, // 2   ******
        8'b11111111, // 3  ********
        8'b11111111, // 4  ********
        8'b01111110, // 5   ******
        8'b00011000, // 6     **
        8'b00000000, // 7
		  // CODE 0x02 - EMPTY BODY ("HALF")
        8'b00000000, // 0
        8'b00011000, // 1     **  
        8'b01111110, // 2   ******
        8'b10000001, // 3  *      *
        8'b10000001, // 4  *      *
        8'b01111110, // 5   ******
        8'b00011000, // 6     **
        8'b00000000, // 7
		  // CODE 0x03 - WHOLE BODY LEFT ("WHOLE")
        8'b00000111, // 0      ***
        8'b00011001, // 1    **  *
        8'b00111000, // 2   ***
        8'b00111000, // 3   ***      
        8'b00111000, // 4   ***      
        8'b00111100, // 5   ****
        8'b00011111, // 6    *****
        8'b00000111, // 7      ***
		  // CODE 0x04 - WHOLE BODY RIGHT ("WHOLE")
        8'b11100000, // 0  ***
        8'b11111000, // 1  *****
        8'b01111100, // 2   *****
        8'b00111100, // 3    ****      
        8'b00111100, // 4    ****      
        8'b00011100, // 5     ***
        8'b00011000, // 6     **
        8'b11100000, // 7  ***
		  // CODE 0x05 - EIGHTH REST TOP
        8'b01000001, // 0   *     *
        8'b11100011, // 1  ***   **
        8'b11100101, // 2  ***  * *
        8'b01111001, // 3   ****  *
        8'b00000010, // 4        *      
        8'b00000010, // 5        *
        8'b00000100, // 6       *
        8'b00000100, // 7       *
		  // CODE 0x06 - EIGHTH REST BOTTOM
        8'b00001000, // 0    *
        8'b00001000, // 1    *
        8'b00010000, // 2   * 
        8'b00010000, // 3   *
        8'b00100000, // 4  *
        8'b00000000, // 5   
        8'b00000000, // 6   
        8'b00000000, // 7    
		  // CODE 0x07 -- QUARTER REST TOP
        8'b00100000, // 0    *
        8'b00010000, // 1     *
        8'b00011000, // 2     **
        8'b00001100, // 3      **  
        8'b00001100, // 4      **   
        8'b00001110, // 5      ***
        8'b00011100, // 6     ***
        8'b00111000, // 7    ***
		  // CODE 0x08 -- QUARTER REST BOTTOM
        8'b00011000, // 0     **
        8'b00001100, // 1      **
        8'b00000110, // 2       **
        8'b00001111, // 3      ****
        8'b00011100, // 4     ***   
        8'b00011000, // 5     **   
        8'b00011000, // 6     **
        8'b00000100, // 7       *
		  // CODE 0x09 - HALF REST LEFT
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00001111, // 2      ****
        8'b00001111, // 3      ****
        8'b00001111, // 4      ****
        8'b00111111, // 5    ******
        8'b00000000, // 6
        8'b00000000, // 7
		  // CODE 0x0A - HALF REST RIGHT
        8'b00000000, // 0
        8'b00000000, // 1
        8'b11110000, // 2  ****
        8'b11110000, // 3  ****
        8'b11110000, // 4  ****
        8'b11111100, // 5  ******
        8'b00000000, // 6
        8'b00000000, // 7
		  // CODE 0x0B - WHOLE REST LEFT
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00111111, // 2    ******
        8'b00001111, // 3      ****
        8'b00001111, // 4      ****
        8'b00001111, // 5      ****
        8'b00000000, // 6
        8'b00000000, // 7
		  // CODE 0x0C - WHOLE REST RIGHT
        8'b00000000, // 0
        8'b00000000, // 1
        8'b11111100, // 2  ******
        8'b11110000, // 3  ****
        8'b11110000, // 4  ****
        8'b11110000, // 5  ****
        8'b00000000, // 6
        8'b00000000, // 7
		  // CODE 0x0D - RESV
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00000000, // 5
        8'b00000000, // 6
        8'b00000000, // 7
		  // CODE 0x0E - RESV
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00000000, // 5
        8'b00000000, // 6
        8'b00000000, // 7
		  // CODE 0x0F - RESV
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00000000, // 5
        8'b00000000, // 6
        8'b00000000, // 7
		  // CODE 0x10 - UP EIGHTH TAIL TOP
        8'b10000000, // 0  *
        8'b10000000, // 1  *
        8'b11000000, // 2  **
        8'b11000000, // 3  **
        8'b11100000, // 4  ***
        8'b11110000, // 5  ****
        8'b00110000, // 6    **
        8'b00011000, // 7     **
		  // CODE 0x11 - UP EIGHTH TAIL BOTTOM
        8'b00001000, // 0      *
        8'b00001000, // 1      *
        8'b00001000, // 2      *
        8'b00001000, // 3      *
        8'b00010000, // 4     *
        8'b00010000, // 5     *
        8'b00100000, // 6    *
        8'b00000000, // 7
		  // CODE 0x12 - DOWN EIGHTH TAIL TOP
        8'b00000000, // 0
        8'b00000100, // 1       *
        8'b00001000, // 2      *
        8'b00001000, // 3      *
        8'b00010000, // 4     *
        8'b00010000, // 5     *
        8'b00010000, // 6     *
        8'b00010000, // 7     *
		  // CODE 0x13 - DOWN EIGHTH TAIL BOTTOM
        8'b00011000, // 0     **
        8'b00001100, // 1      **
        8'b00001111, // 2      ****
        8'b00000111, // 3       ***
        8'b00000011, // 4        **
        8'b00000011, // 5        **
        8'b00000001, // 6         *
        8'b00000001, // 7         *
		  // CODE 0x14 - UP SIXTEENTH TAIL TOP
        8'b10000000, // 0
        8'b11000000, // 1
        8'b01100000, // 2
        8'b10110000, // 3
        8'b11001000, // 4
        8'b00110100, // 5
        8'b00001100, // 6
        8'b00000110, // 7
		  // CODE 0x15 - UP SIXTEENTH TAIL BOTTOM
        8'b00000110, // 0
        8'b00000010, // 1
        8'b00000010, // 2
        8'b00000010, // 3
        8'b00000100, // 4
        8'b00000100, // 5
        8'b00001000, // 6
        8'b00000000, // 7
		  // CODE 0x16 - DOWN SIXTEENTH TAIL TOP
        8'b00000000, // 0
        8'b00010000, // 1
        8'b00100000, // 2
        8'b00100000, // 3
        8'b01000000, // 4
        8'b01000000, // 5
        8'b01000000, // 6
        8'b01100000, // 7
		  // CODE 0x17 - DOWN SIXTEENTH TAIL BOTTOM
        8'b01100000, // 0
        8'b00110000, // 1
        8'b00101100, // 2
        8'b00010011, // 3
        8'b00001101, // 4
        8'b00000110, // 5
        8'b00000011, // 6
        8'b00000001, // 7
		  // CODE 0x18 - SHARP TOP
        8'b00000000, // 0
        8'b00000100, // 1
        8'b00100110, // 2
        8'b00101110, // 3
        8'b00111100, // 4
        8'b00111100, // 5
        8'b01110100, // 6
        8'b01100100, // 7
		  // CODE 0x19 - SHARP BOTTOM
        8'b00100110, // 0
        8'b00101110, // 1
        8'b00111100, // 2
        8'b00111100, // 3
        8'b01110100, // 4
        8'b01100000, // 5
        8'b00100000, // 6
        8'b00000000, // 7
		  // CODE 0x1A - RESV
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00000000, // 5
        8'b00000000, // 6
        8'b00000000, // 7
		  // CODE 0x1B - RESV
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00000000, // 5
        8'b00000000, // 6
        8'b00000000, // 7
		  // CODE 0x1C - RESV
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00000000, // 5
        8'b00000000, // 6
        8'b00000000, // 7
		  // CODE 0x1D - RESV
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00000000, // 5
        8'b00000000, // 6
        8'b00000000, // 7
		  // CODE 0x1E - RESV
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00000000, // 5
        8'b00000000, // 6
        8'b00000000, // 7
		  // CODE 0x1F - RESV
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00000000, // 5
        8'b00000000, // 6
        8'b00000000 // 7
	};
	
	
	assign data = ROM[addr];

endmodule
