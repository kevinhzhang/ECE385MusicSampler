module MusicSampler();
endmodule
